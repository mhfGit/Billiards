library verilog;
use verilog.vl_types.all;
entity blitter is
    port(
        clk             : in     vl_logic;
        reset           : in     vl_logic;
        run             : in     vl_logic;
        oneballx        : in     vl_logic_vector(9 downto 0);
        onebally        : in     vl_logic_vector(9 downto 0);
        twoballx        : in     vl_logic_vector(9 downto 0);
        twobally        : in     vl_logic_vector(9 downto 0);
        threeballx      : in     vl_logic_vector(9 downto 0);
        threebally      : in     vl_logic_vector(9 downto 0);
        fourballx       : in     vl_logic_vector(9 downto 0);
        fourbally       : in     vl_logic_vector(9 downto 0);
        fiveballx       : in     vl_logic_vector(9 downto 0);
        fivebally       : in     vl_logic_vector(9 downto 0);
        sixballx        : in     vl_logic_vector(9 downto 0);
        sixbally        : in     vl_logic_vector(9 downto 0);
        sevenballx      : in     vl_logic_vector(9 downto 0);
        sevenbally      : in     vl_logic_vector(9 downto 0);
        eightballx      : in     vl_logic_vector(9 downto 0);
        eightbally      : in     vl_logic_vector(9 downto 0);
        nineballx       : in     vl_logic_vector(9 downto 0);
        ninebally       : in     vl_logic_vector(9 downto 0);
        tenballx        : in     vl_logic_vector(9 downto 0);
        tenbally        : in     vl_logic_vector(9 downto 0);
        elevenballx     : in     vl_logic_vector(9 downto 0);
        elevenbally     : in     vl_logic_vector(9 downto 0);
        twelveballx     : in     vl_logic_vector(9 downto 0);
        twelvebally     : in     vl_logic_vector(9 downto 0);
        thirteenballx   : in     vl_logic_vector(9 downto 0);
        thirteenbally   : in     vl_logic_vector(9 downto 0);
        fourteenballx   : in     vl_logic_vector(9 downto 0);
        fourteenbally   : in     vl_logic_vector(9 downto 0);
        fifteenballx    : in     vl_logic_vector(9 downto 0);
        fifteenbally    : in     vl_logic_vector(9 downto 0);
        cueballx        : in     vl_logic_vector(9 downto 0);
        cuebally        : in     vl_logic_vector(9 downto 0);
        p1cuex          : in     vl_logic_vector(9 downto 0);
        p1cuey          : in     vl_logic_vector(9 downto 0);
        curpixX         : in     vl_logic_vector(9 downto 0);
        curpixY         : in     vl_logic_vector(9 downto 0);
        direction       : in     vl_logic_vector(2 downto 0);
        to_sw_sig       : out    vl_logic;
        \select\        : out    vl_logic_vector(4 downto 0);
        addrp1cue       : out    vl_logic_vector(15 downto 0);
        addrp1cue45     : out    vl_logic_vector(15 downto 0);
        addrp1cue90     : out    vl_logic_vector(15 downto 0);
        addrp1cue135    : out    vl_logic_vector(15 downto 0);
        addrp1cue180    : out    vl_logic_vector(15 downto 0);
        addrp1cue225    : out    vl_logic_vector(15 downto 0);
        addrp1cue270    : out    vl_logic_vector(15 downto 0);
        addrp1cue315    : out    vl_logic_vector(15 downto 0);
        addrpt          : out    vl_logic_vector(18 downto 0);
        addr1           : out    vl_logic_vector(7 downto 0);
        addr2           : out    vl_logic_vector(7 downto 0);
        addr3           : out    vl_logic_vector(7 downto 0);
        addr4           : out    vl_logic_vector(7 downto 0);
        addr5           : out    vl_logic_vector(7 downto 0);
        addr6           : out    vl_logic_vector(7 downto 0);
        addr7           : out    vl_logic_vector(7 downto 0);
        addr8           : out    vl_logic_vector(7 downto 0);
        addr9           : out    vl_logic_vector(7 downto 0);
        addr10          : out    vl_logic_vector(7 downto 0);
        addr11          : out    vl_logic_vector(7 downto 0);
        addr12          : out    vl_logic_vector(7 downto 0);
        addr13          : out    vl_logic_vector(7 downto 0);
        addr14          : out    vl_logic_vector(7 downto 0);
        addr15          : out    vl_logic_vector(7 downto 0);
        addrcue         : out    vl_logic_vector(7 downto 0);
        collision       : out    vl_logic_vector(16 downto 0)
    );
end blitter;
