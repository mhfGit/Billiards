// nios_system.v

// Generated using ACDS version 14.0 200 at 2015.12.05.22:35:54

`timescale 1 ps / 1 ps
module nios_system (
		input  wire        clk_clk,                //             clk.clk
		output wire [19:0] cueball_export,         //         cueball.export
		output wire [19:0] eightball_export,       //       eightball.export
		output wire [19:0] elevenball_export,      //      elevenball.export
		output wire [19:0] fifteenball_export,     //     fifteenball.export
		output wire [19:0] fiveball_export,        //        fiveball.export
		output wire [19:0] fourball_export,        //        fourball.export
		output wire [19:0] fourteenball_export,    //    fourteenball.export
		output wire [15:0] keycode_export,         //         keycode.export
		output wire [19:0] nineball_export,        //        nineball.export
		output wire [19:0] oneball_export,         //         oneball.export
		output wire [1:0]  otg_hpi_address_export, // otg_hpi_address.export
		output wire        otg_hpi_cs_export,      //      otg_hpi_cs.export
		input  wire [15:0] otg_hpi_data_in_port,   //    otg_hpi_data.in_port
		output wire [15:0] otg_hpi_data_out_port,  //                .out_port
		output wire        otg_hpi_r_export,       //       otg_hpi_r.export
		output wire        otg_hpi_w_export,       //       otg_hpi_w.export
		output wire [19:0] poolcue_export,         //         poolcue.export
		input  wire        reset_reset_n,          //           reset.reset_n
		output wire        sdram_clk_clk,          //       sdram_clk.clk
		output wire [12:0] sdram_wire_addr,        //      sdram_wire.addr
		output wire [1:0]  sdram_wire_ba,          //                .ba
		output wire        sdram_wire_cas_n,       //                .cas_n
		output wire        sdram_wire_cke,         //                .cke
		output wire        sdram_wire_cs_n,        //                .cs_n
		inout  wire [31:0] sdram_wire_dq,          //                .dq
		output wire [3:0]  sdram_wire_dqm,         //                .dqm
		output wire        sdram_wire_ras_n,       //                .ras_n
		output wire        sdram_wire_we_n,        //                .we_n
		output wire [19:0] sevenball_export,       //       sevenball.export
		output wire [19:0] sixball_export,         //         sixball.export
		output wire [19:0] tenball_export,         //         tenball.export
		output wire [19:0] thirteenball_export,    //    thirteenball.export
		output wire [19:0] threeball_export,       //       threeball.export
		output wire [19:0] twelveball_export,      //      twelveball.export
		output wire [19:0] twoball_export,         //         twoball.export
		input  wire        sys_reset_export,       //       sys_reset.export
		input  wire        hw_sig_export,          //          hw_sig.export
		output wire [2:0]  stick_direction_export  // stick_direction.export
	);

	wire         sdram_pll_c0_clk;                                             // sdram_pll:c0 -> [mm_interconnect_0:sdram_pll_c0_clk, rst_controller_002:clk, sdram:clk]
	wire         nios2_qsys_0_data_master_waitrequest;                         // mm_interconnect_0:nios2_qsys_0_data_master_waitrequest -> nios2_qsys_0:d_waitrequest
	wire  [31:0] nios2_qsys_0_data_master_writedata;                           // nios2_qsys_0:d_writedata -> mm_interconnect_0:nios2_qsys_0_data_master_writedata
	wire  [28:0] nios2_qsys_0_data_master_address;                             // nios2_qsys_0:d_address -> mm_interconnect_0:nios2_qsys_0_data_master_address
	wire         nios2_qsys_0_data_master_write;                               // nios2_qsys_0:d_write -> mm_interconnect_0:nios2_qsys_0_data_master_write
	wire         nios2_qsys_0_data_master_read;                                // nios2_qsys_0:d_read -> mm_interconnect_0:nios2_qsys_0_data_master_read
	wire  [31:0] nios2_qsys_0_data_master_readdata;                            // mm_interconnect_0:nios2_qsys_0_data_master_readdata -> nios2_qsys_0:d_readdata
	wire         nios2_qsys_0_data_master_debugaccess;                         // nios2_qsys_0:jtag_debug_module_debugaccess_to_roms -> mm_interconnect_0:nios2_qsys_0_data_master_debugaccess
	wire   [3:0] nios2_qsys_0_data_master_byteenable;                          // nios2_qsys_0:d_byteenable -> mm_interconnect_0:nios2_qsys_0_data_master_byteenable
	wire         nios2_qsys_0_instruction_master_waitrequest;                  // mm_interconnect_0:nios2_qsys_0_instruction_master_waitrequest -> nios2_qsys_0:i_waitrequest
	wire  [28:0] nios2_qsys_0_instruction_master_address;                      // nios2_qsys_0:i_address -> mm_interconnect_0:nios2_qsys_0_instruction_master_address
	wire         nios2_qsys_0_instruction_master_read;                         // nios2_qsys_0:i_read -> mm_interconnect_0:nios2_qsys_0_instruction_master_read
	wire  [31:0] nios2_qsys_0_instruction_master_readdata;                     // mm_interconnect_0:nios2_qsys_0_instruction_master_readdata -> nios2_qsys_0:i_readdata
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest;  // jtag_uart_0:av_waitrequest -> mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_waitrequest
	wire  [31:0] mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata;    // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_writedata -> jtag_uart_0:av_writedata
	wire   [0:0] mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address;      // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_address -> jtag_uart_0:av_address
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect;   // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_chipselect -> jtag_uart_0:av_chipselect
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write;        // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_write -> jtag_uart_0:av_write_n
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read;         // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_read -> jtag_uart_0:av_read_n
	wire  [31:0] mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata;     // jtag_uart_0:av_readdata -> mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_readdata
	wire   [0:0] mm_interconnect_0_sysid_qsys_0_control_slave_address;         // mm_interconnect_0:sysid_qsys_0_control_slave_address -> sysid_qsys_0:address
	wire  [31:0] mm_interconnect_0_sysid_qsys_0_control_slave_readdata;        // sysid_qsys_0:readdata -> mm_interconnect_0:sysid_qsys_0_control_slave_readdata
	wire         mm_interconnect_0_nios2_qsys_0_jtag_debug_module_waitrequest; // nios2_qsys_0:jtag_debug_module_waitrequest -> mm_interconnect_0:nios2_qsys_0_jtag_debug_module_waitrequest
	wire  [31:0] mm_interconnect_0_nios2_qsys_0_jtag_debug_module_writedata;   // mm_interconnect_0:nios2_qsys_0_jtag_debug_module_writedata -> nios2_qsys_0:jtag_debug_module_writedata
	wire   [8:0] mm_interconnect_0_nios2_qsys_0_jtag_debug_module_address;     // mm_interconnect_0:nios2_qsys_0_jtag_debug_module_address -> nios2_qsys_0:jtag_debug_module_address
	wire         mm_interconnect_0_nios2_qsys_0_jtag_debug_module_write;       // mm_interconnect_0:nios2_qsys_0_jtag_debug_module_write -> nios2_qsys_0:jtag_debug_module_write
	wire         mm_interconnect_0_nios2_qsys_0_jtag_debug_module_read;        // mm_interconnect_0:nios2_qsys_0_jtag_debug_module_read -> nios2_qsys_0:jtag_debug_module_read
	wire  [31:0] mm_interconnect_0_nios2_qsys_0_jtag_debug_module_readdata;    // nios2_qsys_0:jtag_debug_module_readdata -> mm_interconnect_0:nios2_qsys_0_jtag_debug_module_readdata
	wire         mm_interconnect_0_nios2_qsys_0_jtag_debug_module_debugaccess; // mm_interconnect_0:nios2_qsys_0_jtag_debug_module_debugaccess -> nios2_qsys_0:jtag_debug_module_debugaccess
	wire   [3:0] mm_interconnect_0_nios2_qsys_0_jtag_debug_module_byteenable;  // mm_interconnect_0:nios2_qsys_0_jtag_debug_module_byteenable -> nios2_qsys_0:jtag_debug_module_byteenable
	wire  [31:0] mm_interconnect_0_sdram_pll_pll_slave_writedata;              // mm_interconnect_0:sdram_pll_pll_slave_writedata -> sdram_pll:writedata
	wire   [1:0] mm_interconnect_0_sdram_pll_pll_slave_address;                // mm_interconnect_0:sdram_pll_pll_slave_address -> sdram_pll:address
	wire         mm_interconnect_0_sdram_pll_pll_slave_write;                  // mm_interconnect_0:sdram_pll_pll_slave_write -> sdram_pll:write
	wire         mm_interconnect_0_sdram_pll_pll_slave_read;                   // mm_interconnect_0:sdram_pll_pll_slave_read -> sdram_pll:read
	wire  [31:0] mm_interconnect_0_sdram_pll_pll_slave_readdata;               // sdram_pll:readdata -> mm_interconnect_0:sdram_pll_pll_slave_readdata
	wire  [31:0] mm_interconnect_0_onchip_memory2_0_s1_writedata;              // mm_interconnect_0:onchip_memory2_0_s1_writedata -> onchip_memory2_0:writedata
	wire   [1:0] mm_interconnect_0_onchip_memory2_0_s1_address;                // mm_interconnect_0:onchip_memory2_0_s1_address -> onchip_memory2_0:address
	wire         mm_interconnect_0_onchip_memory2_0_s1_chipselect;             // mm_interconnect_0:onchip_memory2_0_s1_chipselect -> onchip_memory2_0:chipselect
	wire         mm_interconnect_0_onchip_memory2_0_s1_clken;                  // mm_interconnect_0:onchip_memory2_0_s1_clken -> onchip_memory2_0:clken
	wire         mm_interconnect_0_onchip_memory2_0_s1_write;                  // mm_interconnect_0:onchip_memory2_0_s1_write -> onchip_memory2_0:write
	wire  [31:0] mm_interconnect_0_onchip_memory2_0_s1_readdata;               // onchip_memory2_0:readdata -> mm_interconnect_0:onchip_memory2_0_s1_readdata
	wire   [3:0] mm_interconnect_0_onchip_memory2_0_s1_byteenable;             // mm_interconnect_0:onchip_memory2_0_s1_byteenable -> onchip_memory2_0:byteenable
	wire         mm_interconnect_0_sdram_s1_waitrequest;                       // sdram:za_waitrequest -> mm_interconnect_0:sdram_s1_waitrequest
	wire  [31:0] mm_interconnect_0_sdram_s1_writedata;                         // mm_interconnect_0:sdram_s1_writedata -> sdram:az_data
	wire  [24:0] mm_interconnect_0_sdram_s1_address;                           // mm_interconnect_0:sdram_s1_address -> sdram:az_addr
	wire         mm_interconnect_0_sdram_s1_chipselect;                        // mm_interconnect_0:sdram_s1_chipselect -> sdram:az_cs
	wire         mm_interconnect_0_sdram_s1_write;                             // mm_interconnect_0:sdram_s1_write -> sdram:az_wr_n
	wire         mm_interconnect_0_sdram_s1_read;                              // mm_interconnect_0:sdram_s1_read -> sdram:az_rd_n
	wire  [31:0] mm_interconnect_0_sdram_s1_readdata;                          // sdram:za_data -> mm_interconnect_0:sdram_s1_readdata
	wire         mm_interconnect_0_sdram_s1_readdatavalid;                     // sdram:za_valid -> mm_interconnect_0:sdram_s1_readdatavalid
	wire   [3:0] mm_interconnect_0_sdram_s1_byteenable;                        // mm_interconnect_0:sdram_s1_byteenable -> sdram:az_be_n
	wire  [31:0] mm_interconnect_0_keycode_s1_writedata;                       // mm_interconnect_0:keycode_s1_writedata -> keycode:writedata
	wire   [1:0] mm_interconnect_0_keycode_s1_address;                         // mm_interconnect_0:keycode_s1_address -> keycode:address
	wire         mm_interconnect_0_keycode_s1_chipselect;                      // mm_interconnect_0:keycode_s1_chipselect -> keycode:chipselect
	wire         mm_interconnect_0_keycode_s1_write;                           // mm_interconnect_0:keycode_s1_write -> keycode:write_n
	wire  [31:0] mm_interconnect_0_keycode_s1_readdata;                        // keycode:readdata -> mm_interconnect_0:keycode_s1_readdata
	wire  [31:0] mm_interconnect_0_otg_hpi_cs_s1_writedata;                    // mm_interconnect_0:otg_hpi_cs_s1_writedata -> otg_hpi_cs:writedata
	wire   [1:0] mm_interconnect_0_otg_hpi_cs_s1_address;                      // mm_interconnect_0:otg_hpi_cs_s1_address -> otg_hpi_cs:address
	wire         mm_interconnect_0_otg_hpi_cs_s1_chipselect;                   // mm_interconnect_0:otg_hpi_cs_s1_chipselect -> otg_hpi_cs:chipselect
	wire         mm_interconnect_0_otg_hpi_cs_s1_write;                        // mm_interconnect_0:otg_hpi_cs_s1_write -> otg_hpi_cs:write_n
	wire  [31:0] mm_interconnect_0_otg_hpi_cs_s1_readdata;                     // otg_hpi_cs:readdata -> mm_interconnect_0:otg_hpi_cs_s1_readdata
	wire  [31:0] mm_interconnect_0_otg_hpi_address_s1_writedata;               // mm_interconnect_0:otg_hpi_address_s1_writedata -> otg_hpi_address:writedata
	wire   [1:0] mm_interconnect_0_otg_hpi_address_s1_address;                 // mm_interconnect_0:otg_hpi_address_s1_address -> otg_hpi_address:address
	wire         mm_interconnect_0_otg_hpi_address_s1_chipselect;              // mm_interconnect_0:otg_hpi_address_s1_chipselect -> otg_hpi_address:chipselect
	wire         mm_interconnect_0_otg_hpi_address_s1_write;                   // mm_interconnect_0:otg_hpi_address_s1_write -> otg_hpi_address:write_n
	wire  [31:0] mm_interconnect_0_otg_hpi_address_s1_readdata;                // otg_hpi_address:readdata -> mm_interconnect_0:otg_hpi_address_s1_readdata
	wire  [31:0] mm_interconnect_0_otg_hpi_data_s1_writedata;                  // mm_interconnect_0:otg_hpi_data_s1_writedata -> otg_hpi_data:writedata
	wire   [1:0] mm_interconnect_0_otg_hpi_data_s1_address;                    // mm_interconnect_0:otg_hpi_data_s1_address -> otg_hpi_data:address
	wire         mm_interconnect_0_otg_hpi_data_s1_chipselect;                 // mm_interconnect_0:otg_hpi_data_s1_chipselect -> otg_hpi_data:chipselect
	wire         mm_interconnect_0_otg_hpi_data_s1_write;                      // mm_interconnect_0:otg_hpi_data_s1_write -> otg_hpi_data:write_n
	wire  [31:0] mm_interconnect_0_otg_hpi_data_s1_readdata;                   // otg_hpi_data:readdata -> mm_interconnect_0:otg_hpi_data_s1_readdata
	wire  [31:0] mm_interconnect_0_otg_hpi_r_s1_writedata;                     // mm_interconnect_0:otg_hpi_r_s1_writedata -> otg_hpi_r:writedata
	wire   [1:0] mm_interconnect_0_otg_hpi_r_s1_address;                       // mm_interconnect_0:otg_hpi_r_s1_address -> otg_hpi_r:address
	wire         mm_interconnect_0_otg_hpi_r_s1_chipselect;                    // mm_interconnect_0:otg_hpi_r_s1_chipselect -> otg_hpi_r:chipselect
	wire         mm_interconnect_0_otg_hpi_r_s1_write;                         // mm_interconnect_0:otg_hpi_r_s1_write -> otg_hpi_r:write_n
	wire  [31:0] mm_interconnect_0_otg_hpi_r_s1_readdata;                      // otg_hpi_r:readdata -> mm_interconnect_0:otg_hpi_r_s1_readdata
	wire  [31:0] mm_interconnect_0_otg_hpi_w_s1_writedata;                     // mm_interconnect_0:otg_hpi_w_s1_writedata -> otg_hpi_w:writedata
	wire   [1:0] mm_interconnect_0_otg_hpi_w_s1_address;                       // mm_interconnect_0:otg_hpi_w_s1_address -> otg_hpi_w:address
	wire         mm_interconnect_0_otg_hpi_w_s1_chipselect;                    // mm_interconnect_0:otg_hpi_w_s1_chipselect -> otg_hpi_w:chipselect
	wire         mm_interconnect_0_otg_hpi_w_s1_write;                         // mm_interconnect_0:otg_hpi_w_s1_write -> otg_hpi_w:write_n
	wire  [31:0] mm_interconnect_0_otg_hpi_w_s1_readdata;                      // otg_hpi_w:readdata -> mm_interconnect_0:otg_hpi_w_s1_readdata
	wire  [31:0] mm_interconnect_0_oneball_s1_writedata;                       // mm_interconnect_0:OneBall_s1_writedata -> OneBall:writedata
	wire   [1:0] mm_interconnect_0_oneball_s1_address;                         // mm_interconnect_0:OneBall_s1_address -> OneBall:address
	wire         mm_interconnect_0_oneball_s1_chipselect;                      // mm_interconnect_0:OneBall_s1_chipselect -> OneBall:chipselect
	wire         mm_interconnect_0_oneball_s1_write;                           // mm_interconnect_0:OneBall_s1_write -> OneBall:write_n
	wire  [31:0] mm_interconnect_0_oneball_s1_readdata;                        // OneBall:readdata -> mm_interconnect_0:OneBall_s1_readdata
	wire  [31:0] mm_interconnect_0_twoball_s1_writedata;                       // mm_interconnect_0:TwoBall_s1_writedata -> TwoBall:writedata
	wire   [1:0] mm_interconnect_0_twoball_s1_address;                         // mm_interconnect_0:TwoBall_s1_address -> TwoBall:address
	wire         mm_interconnect_0_twoball_s1_chipselect;                      // mm_interconnect_0:TwoBall_s1_chipselect -> TwoBall:chipselect
	wire         mm_interconnect_0_twoball_s1_write;                           // mm_interconnect_0:TwoBall_s1_write -> TwoBall:write_n
	wire  [31:0] mm_interconnect_0_twoball_s1_readdata;                        // TwoBall:readdata -> mm_interconnect_0:TwoBall_s1_readdata
	wire  [31:0] mm_interconnect_0_threeball_s1_writedata;                     // mm_interconnect_0:ThreeBall_s1_writedata -> ThreeBall:writedata
	wire   [1:0] mm_interconnect_0_threeball_s1_address;                       // mm_interconnect_0:ThreeBall_s1_address -> ThreeBall:address
	wire         mm_interconnect_0_threeball_s1_chipselect;                    // mm_interconnect_0:ThreeBall_s1_chipselect -> ThreeBall:chipselect
	wire         mm_interconnect_0_threeball_s1_write;                         // mm_interconnect_0:ThreeBall_s1_write -> ThreeBall:write_n
	wire  [31:0] mm_interconnect_0_threeball_s1_readdata;                      // ThreeBall:readdata -> mm_interconnect_0:ThreeBall_s1_readdata
	wire  [31:0] mm_interconnect_0_fourball_s1_writedata;                      // mm_interconnect_0:FourBall_s1_writedata -> FourBall:writedata
	wire   [1:0] mm_interconnect_0_fourball_s1_address;                        // mm_interconnect_0:FourBall_s1_address -> FourBall:address
	wire         mm_interconnect_0_fourball_s1_chipselect;                     // mm_interconnect_0:FourBall_s1_chipselect -> FourBall:chipselect
	wire         mm_interconnect_0_fourball_s1_write;                          // mm_interconnect_0:FourBall_s1_write -> FourBall:write_n
	wire  [31:0] mm_interconnect_0_fourball_s1_readdata;                       // FourBall:readdata -> mm_interconnect_0:FourBall_s1_readdata
	wire  [31:0] mm_interconnect_0_fiveball_s1_writedata;                      // mm_interconnect_0:FiveBall_s1_writedata -> FiveBall:writedata
	wire   [1:0] mm_interconnect_0_fiveball_s1_address;                        // mm_interconnect_0:FiveBall_s1_address -> FiveBall:address
	wire         mm_interconnect_0_fiveball_s1_chipselect;                     // mm_interconnect_0:FiveBall_s1_chipselect -> FiveBall:chipselect
	wire         mm_interconnect_0_fiveball_s1_write;                          // mm_interconnect_0:FiveBall_s1_write -> FiveBall:write_n
	wire  [31:0] mm_interconnect_0_fiveball_s1_readdata;                       // FiveBall:readdata -> mm_interconnect_0:FiveBall_s1_readdata
	wire  [31:0] mm_interconnect_0_sixball_s1_writedata;                       // mm_interconnect_0:SixBall_s1_writedata -> SixBall:writedata
	wire   [1:0] mm_interconnect_0_sixball_s1_address;                         // mm_interconnect_0:SixBall_s1_address -> SixBall:address
	wire         mm_interconnect_0_sixball_s1_chipselect;                      // mm_interconnect_0:SixBall_s1_chipselect -> SixBall:chipselect
	wire         mm_interconnect_0_sixball_s1_write;                           // mm_interconnect_0:SixBall_s1_write -> SixBall:write_n
	wire  [31:0] mm_interconnect_0_sixball_s1_readdata;                        // SixBall:readdata -> mm_interconnect_0:SixBall_s1_readdata
	wire  [31:0] mm_interconnect_0_sevenball_s1_writedata;                     // mm_interconnect_0:SevenBall_s1_writedata -> SevenBall:writedata
	wire   [1:0] mm_interconnect_0_sevenball_s1_address;                       // mm_interconnect_0:SevenBall_s1_address -> SevenBall:address
	wire         mm_interconnect_0_sevenball_s1_chipselect;                    // mm_interconnect_0:SevenBall_s1_chipselect -> SevenBall:chipselect
	wire         mm_interconnect_0_sevenball_s1_write;                         // mm_interconnect_0:SevenBall_s1_write -> SevenBall:write_n
	wire  [31:0] mm_interconnect_0_sevenball_s1_readdata;                      // SevenBall:readdata -> mm_interconnect_0:SevenBall_s1_readdata
	wire  [31:0] mm_interconnect_0_eightball_s1_writedata;                     // mm_interconnect_0:EightBall_s1_writedata -> EightBall:writedata
	wire   [1:0] mm_interconnect_0_eightball_s1_address;                       // mm_interconnect_0:EightBall_s1_address -> EightBall:address
	wire         mm_interconnect_0_eightball_s1_chipselect;                    // mm_interconnect_0:EightBall_s1_chipselect -> EightBall:chipselect
	wire         mm_interconnect_0_eightball_s1_write;                         // mm_interconnect_0:EightBall_s1_write -> EightBall:write_n
	wire  [31:0] mm_interconnect_0_eightball_s1_readdata;                      // EightBall:readdata -> mm_interconnect_0:EightBall_s1_readdata
	wire  [31:0] mm_interconnect_0_nineball_s1_writedata;                      // mm_interconnect_0:NineBall_s1_writedata -> NineBall:writedata
	wire   [1:0] mm_interconnect_0_nineball_s1_address;                        // mm_interconnect_0:NineBall_s1_address -> NineBall:address
	wire         mm_interconnect_0_nineball_s1_chipselect;                     // mm_interconnect_0:NineBall_s1_chipselect -> NineBall:chipselect
	wire         mm_interconnect_0_nineball_s1_write;                          // mm_interconnect_0:NineBall_s1_write -> NineBall:write_n
	wire  [31:0] mm_interconnect_0_nineball_s1_readdata;                       // NineBall:readdata -> mm_interconnect_0:NineBall_s1_readdata
	wire  [31:0] mm_interconnect_0_tenball_s1_writedata;                       // mm_interconnect_0:TenBall_s1_writedata -> TenBall:writedata
	wire   [1:0] mm_interconnect_0_tenball_s1_address;                         // mm_interconnect_0:TenBall_s1_address -> TenBall:address
	wire         mm_interconnect_0_tenball_s1_chipselect;                      // mm_interconnect_0:TenBall_s1_chipselect -> TenBall:chipselect
	wire         mm_interconnect_0_tenball_s1_write;                           // mm_interconnect_0:TenBall_s1_write -> TenBall:write_n
	wire  [31:0] mm_interconnect_0_tenball_s1_readdata;                        // TenBall:readdata -> mm_interconnect_0:TenBall_s1_readdata
	wire  [31:0] mm_interconnect_0_elevenball_s1_writedata;                    // mm_interconnect_0:ElevenBall_s1_writedata -> ElevenBall:writedata
	wire   [1:0] mm_interconnect_0_elevenball_s1_address;                      // mm_interconnect_0:ElevenBall_s1_address -> ElevenBall:address
	wire         mm_interconnect_0_elevenball_s1_chipselect;                   // mm_interconnect_0:ElevenBall_s1_chipselect -> ElevenBall:chipselect
	wire         mm_interconnect_0_elevenball_s1_write;                        // mm_interconnect_0:ElevenBall_s1_write -> ElevenBall:write_n
	wire  [31:0] mm_interconnect_0_elevenball_s1_readdata;                     // ElevenBall:readdata -> mm_interconnect_0:ElevenBall_s1_readdata
	wire  [31:0] mm_interconnect_0_twelveball_s1_writedata;                    // mm_interconnect_0:TwelveBall_s1_writedata -> TwelveBall:writedata
	wire   [1:0] mm_interconnect_0_twelveball_s1_address;                      // mm_interconnect_0:TwelveBall_s1_address -> TwelveBall:address
	wire         mm_interconnect_0_twelveball_s1_chipselect;                   // mm_interconnect_0:TwelveBall_s1_chipselect -> TwelveBall:chipselect
	wire         mm_interconnect_0_twelveball_s1_write;                        // mm_interconnect_0:TwelveBall_s1_write -> TwelveBall:write_n
	wire  [31:0] mm_interconnect_0_twelveball_s1_readdata;                     // TwelveBall:readdata -> mm_interconnect_0:TwelveBall_s1_readdata
	wire  [31:0] mm_interconnect_0_thirteenball_s1_writedata;                  // mm_interconnect_0:ThirteenBall_s1_writedata -> ThirteenBall:writedata
	wire   [1:0] mm_interconnect_0_thirteenball_s1_address;                    // mm_interconnect_0:ThirteenBall_s1_address -> ThirteenBall:address
	wire         mm_interconnect_0_thirteenball_s1_chipselect;                 // mm_interconnect_0:ThirteenBall_s1_chipselect -> ThirteenBall:chipselect
	wire         mm_interconnect_0_thirteenball_s1_write;                      // mm_interconnect_0:ThirteenBall_s1_write -> ThirteenBall:write_n
	wire  [31:0] mm_interconnect_0_thirteenball_s1_readdata;                   // ThirteenBall:readdata -> mm_interconnect_0:ThirteenBall_s1_readdata
	wire  [31:0] mm_interconnect_0_fourteenball_s1_writedata;                  // mm_interconnect_0:FourteenBall_s1_writedata -> FourteenBall:writedata
	wire   [1:0] mm_interconnect_0_fourteenball_s1_address;                    // mm_interconnect_0:FourteenBall_s1_address -> FourteenBall:address
	wire         mm_interconnect_0_fourteenball_s1_chipselect;                 // mm_interconnect_0:FourteenBall_s1_chipselect -> FourteenBall:chipselect
	wire         mm_interconnect_0_fourteenball_s1_write;                      // mm_interconnect_0:FourteenBall_s1_write -> FourteenBall:write_n
	wire  [31:0] mm_interconnect_0_fourteenball_s1_readdata;                   // FourteenBall:readdata -> mm_interconnect_0:FourteenBall_s1_readdata
	wire  [31:0] mm_interconnect_0_fifteenball_s1_writedata;                   // mm_interconnect_0:FifteenBall_s1_writedata -> FifteenBall:writedata
	wire   [1:0] mm_interconnect_0_fifteenball_s1_address;                     // mm_interconnect_0:FifteenBall_s1_address -> FifteenBall:address
	wire         mm_interconnect_0_fifteenball_s1_chipselect;                  // mm_interconnect_0:FifteenBall_s1_chipselect -> FifteenBall:chipselect
	wire         mm_interconnect_0_fifteenball_s1_write;                       // mm_interconnect_0:FifteenBall_s1_write -> FifteenBall:write_n
	wire  [31:0] mm_interconnect_0_fifteenball_s1_readdata;                    // FifteenBall:readdata -> mm_interconnect_0:FifteenBall_s1_readdata
	wire  [31:0] mm_interconnect_0_cueball_s1_writedata;                       // mm_interconnect_0:cueBall_s1_writedata -> cueBall:writedata
	wire   [1:0] mm_interconnect_0_cueball_s1_address;                         // mm_interconnect_0:cueBall_s1_address -> cueBall:address
	wire         mm_interconnect_0_cueball_s1_chipselect;                      // mm_interconnect_0:cueBall_s1_chipselect -> cueBall:chipselect
	wire         mm_interconnect_0_cueball_s1_write;                           // mm_interconnect_0:cueBall_s1_write -> cueBall:write_n
	wire  [31:0] mm_interconnect_0_cueball_s1_readdata;                        // cueBall:readdata -> mm_interconnect_0:cueBall_s1_readdata
	wire  [31:0] mm_interconnect_0_poolcue_s1_writedata;                       // mm_interconnect_0:poolcue_s1_writedata -> poolcue:writedata
	wire   [1:0] mm_interconnect_0_poolcue_s1_address;                         // mm_interconnect_0:poolcue_s1_address -> poolcue:address
	wire         mm_interconnect_0_poolcue_s1_chipselect;                      // mm_interconnect_0:poolcue_s1_chipselect -> poolcue:chipselect
	wire         mm_interconnect_0_poolcue_s1_write;                           // mm_interconnect_0:poolcue_s1_write -> poolcue:write_n
	wire  [31:0] mm_interconnect_0_poolcue_s1_readdata;                        // poolcue:readdata -> mm_interconnect_0:poolcue_s1_readdata
	wire   [1:0] mm_interconnect_0_reset_s1_address;                           // mm_interconnect_0:reset_s1_address -> reset:address
	wire  [31:0] mm_interconnect_0_reset_s1_readdata;                          // reset:readdata -> mm_interconnect_0:reset_s1_readdata
	wire   [1:0] mm_interconnect_0_hw_sig_s1_address;                          // mm_interconnect_0:hw_sig_s1_address -> hw_sig:address
	wire  [31:0] mm_interconnect_0_hw_sig_s1_readdata;                         // hw_sig:readdata -> mm_interconnect_0:hw_sig_s1_readdata
	wire  [31:0] mm_interconnect_0_stick_direction_s1_writedata;               // mm_interconnect_0:stick_direction_s1_writedata -> stick_direction:writedata
	wire   [1:0] mm_interconnect_0_stick_direction_s1_address;                 // mm_interconnect_0:stick_direction_s1_address -> stick_direction:address
	wire         mm_interconnect_0_stick_direction_s1_chipselect;              // mm_interconnect_0:stick_direction_s1_chipselect -> stick_direction:chipselect
	wire         mm_interconnect_0_stick_direction_s1_write;                   // mm_interconnect_0:stick_direction_s1_write -> stick_direction:write_n
	wire  [31:0] mm_interconnect_0_stick_direction_s1_readdata;                // stick_direction:readdata -> mm_interconnect_0:stick_direction_s1_readdata
	wire         irq_mapper_receiver0_irq;                                     // jtag_uart_0:av_irq -> irq_mapper:receiver0_irq
	wire  [31:0] nios2_qsys_0_d_irq_irq;                                       // irq_mapper:sender_irq -> nios2_qsys_0:d_irq
	wire         rst_controller_reset_out_reset;                               // rst_controller:reset_out -> [EightBall:reset_n, ElevenBall:reset_n, FifteenBall:reset_n, FiveBall:reset_n, FourBall:reset_n, FourteenBall:reset_n, NineBall:reset_n, OneBall:reset_n, SevenBall:reset_n, SixBall:reset_n, TenBall:reset_n, ThirteenBall:reset_n, ThreeBall:reset_n, TwelveBall:reset_n, TwoBall:reset_n, cueBall:reset_n, hw_sig:reset_n, jtag_uart_0:rst_n, keycode:reset_n, mm_interconnect_0:jtag_uart_0_reset_reset_bridge_in_reset_reset, otg_hpi_address:reset_n, otg_hpi_cs:reset_n, otg_hpi_data:reset_n, otg_hpi_r:reset_n, otg_hpi_w:reset_n, poolcue:reset_n, reset:reset_n, stick_direction:reset_n]
	wire         nios2_qsys_0_jtag_debug_module_reset_reset;                   // nios2_qsys_0:jtag_debug_module_resetrequest -> rst_controller:reset_in1
	wire         rst_controller_001_reset_out_reset;                           // rst_controller_001:reset_out -> [irq_mapper:reset, mm_interconnect_0:nios2_qsys_0_reset_n_reset_bridge_in_reset_reset, nios2_qsys_0:reset_n, onchip_memory2_0:reset, rst_translator:in_reset, sdram_pll:reset, sysid_qsys_0:reset_n]
	wire         rst_controller_001_reset_out_reset_req;                       // rst_controller_001:reset_req -> [nios2_qsys_0:reset_req, onchip_memory2_0:reset_req, rst_translator:reset_req_in]
	wire         rst_controller_002_reset_out_reset;                           // rst_controller_002:reset_out -> [mm_interconnect_0:sdram_reset_reset_bridge_in_reset_reset, sdram:reset_n]

	nios_system_EightBall eightball (
		.clk        (clk_clk),                                   //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),           //               reset.reset_n
		.address    (mm_interconnect_0_eightball_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_eightball_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_eightball_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_eightball_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_eightball_s1_readdata),   //                    .readdata
		.out_port   (eightball_export)                           // external_connection.export
	);

	nios_system_EightBall elevenball (
		.clk        (clk_clk),                                    //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),            //               reset.reset_n
		.address    (mm_interconnect_0_elevenball_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_elevenball_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_elevenball_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_elevenball_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_elevenball_s1_readdata),   //                    .readdata
		.out_port   (elevenball_export)                           // external_connection.export
	);

	nios_system_EightBall fifteenball (
		.clk        (clk_clk),                                     //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),             //               reset.reset_n
		.address    (mm_interconnect_0_fifteenball_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_fifteenball_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_fifteenball_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_fifteenball_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_fifteenball_s1_readdata),   //                    .readdata
		.out_port   (fifteenball_export)                           // external_connection.export
	);

	nios_system_EightBall fiveball (
		.clk        (clk_clk),                                  //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),          //               reset.reset_n
		.address    (mm_interconnect_0_fiveball_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_fiveball_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_fiveball_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_fiveball_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_fiveball_s1_readdata),   //                    .readdata
		.out_port   (fiveball_export)                           // external_connection.export
	);

	nios_system_EightBall fourball (
		.clk        (clk_clk),                                  //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),          //               reset.reset_n
		.address    (mm_interconnect_0_fourball_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_fourball_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_fourball_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_fourball_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_fourball_s1_readdata),   //                    .readdata
		.out_port   (fourball_export)                           // external_connection.export
	);

	nios_system_EightBall fourteenball (
		.clk        (clk_clk),                                      //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),              //               reset.reset_n
		.address    (mm_interconnect_0_fourteenball_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_fourteenball_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_fourteenball_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_fourteenball_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_fourteenball_s1_readdata),   //                    .readdata
		.out_port   (fourteenball_export)                           // external_connection.export
	);

	nios_system_EightBall nineball (
		.clk        (clk_clk),                                  //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),          //               reset.reset_n
		.address    (mm_interconnect_0_nineball_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_nineball_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_nineball_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_nineball_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_nineball_s1_readdata),   //                    .readdata
		.out_port   (nineball_export)                           // external_connection.export
	);

	nios_system_EightBall oneball (
		.clk        (clk_clk),                                 //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),         //               reset.reset_n
		.address    (mm_interconnect_0_oneball_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_oneball_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_oneball_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_oneball_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_oneball_s1_readdata),   //                    .readdata
		.out_port   (oneball_export)                           // external_connection.export
	);

	nios_system_EightBall sevenball (
		.clk        (clk_clk),                                   //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),           //               reset.reset_n
		.address    (mm_interconnect_0_sevenball_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_sevenball_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_sevenball_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_sevenball_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_sevenball_s1_readdata),   //                    .readdata
		.out_port   (sevenball_export)                           // external_connection.export
	);

	nios_system_EightBall sixball (
		.clk        (clk_clk),                                 //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),         //               reset.reset_n
		.address    (mm_interconnect_0_sixball_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_sixball_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_sixball_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_sixball_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_sixball_s1_readdata),   //                    .readdata
		.out_port   (sixball_export)                           // external_connection.export
	);

	nios_system_EightBall tenball (
		.clk        (clk_clk),                                 //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),         //               reset.reset_n
		.address    (mm_interconnect_0_tenball_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_tenball_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_tenball_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_tenball_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_tenball_s1_readdata),   //                    .readdata
		.out_port   (tenball_export)                           // external_connection.export
	);

	nios_system_EightBall thirteenball (
		.clk        (clk_clk),                                      //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),              //               reset.reset_n
		.address    (mm_interconnect_0_thirteenball_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_thirteenball_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_thirteenball_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_thirteenball_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_thirteenball_s1_readdata),   //                    .readdata
		.out_port   (thirteenball_export)                           // external_connection.export
	);

	nios_system_EightBall threeball (
		.clk        (clk_clk),                                   //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),           //               reset.reset_n
		.address    (mm_interconnect_0_threeball_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_threeball_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_threeball_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_threeball_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_threeball_s1_readdata),   //                    .readdata
		.out_port   (threeball_export)                           // external_connection.export
	);

	nios_system_EightBall twelveball (
		.clk        (clk_clk),                                    //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),            //               reset.reset_n
		.address    (mm_interconnect_0_twelveball_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_twelveball_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_twelveball_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_twelveball_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_twelveball_s1_readdata),   //                    .readdata
		.out_port   (twelveball_export)                           // external_connection.export
	);

	nios_system_EightBall twoball (
		.clk        (clk_clk),                                 //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),         //               reset.reset_n
		.address    (mm_interconnect_0_twoball_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_twoball_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_twoball_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_twoball_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_twoball_s1_readdata),   //                    .readdata
		.out_port   (twoball_export)                           // external_connection.export
	);

	nios_system_EightBall cueball (
		.clk        (clk_clk),                                 //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),         //               reset.reset_n
		.address    (mm_interconnect_0_cueball_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_cueball_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_cueball_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_cueball_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_cueball_s1_readdata),   //                    .readdata
		.out_port   (cueball_export)                           // external_connection.export
	);

	nios_system_jtag_uart_0 jtag_uart_0 (
		.clk            (clk_clk),                                                     //               clk.clk
		.rst_n          (~rst_controller_reset_out_reset),                             //             reset.reset_n
		.av_chipselect  (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver0_irq)                                     //               irq.irq
	);

	nios_system_keycode keycode (
		.clk        (clk_clk),                                 //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),         //               reset.reset_n
		.address    (mm_interconnect_0_keycode_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_keycode_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_keycode_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_keycode_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_keycode_s1_readdata),   //                    .readdata
		.out_port   (keycode_export)                           // external_connection.export
	);

	nios_system_nios2_qsys_0 nios2_qsys_0 (
		.clk                                   (clk_clk),                                                      //                       clk.clk
		.reset_n                               (~rst_controller_001_reset_out_reset),                          //                   reset_n.reset_n
		.reset_req                             (rst_controller_001_reset_out_reset_req),                       //                          .reset_req
		.d_address                             (nios2_qsys_0_data_master_address),                             //               data_master.address
		.d_byteenable                          (nios2_qsys_0_data_master_byteenable),                          //                          .byteenable
		.d_read                                (nios2_qsys_0_data_master_read),                                //                          .read
		.d_readdata                            (nios2_qsys_0_data_master_readdata),                            //                          .readdata
		.d_waitrequest                         (nios2_qsys_0_data_master_waitrequest),                         //                          .waitrequest
		.d_write                               (nios2_qsys_0_data_master_write),                               //                          .write
		.d_writedata                           (nios2_qsys_0_data_master_writedata),                           //                          .writedata
		.jtag_debug_module_debugaccess_to_roms (nios2_qsys_0_data_master_debugaccess),                         //                          .debugaccess
		.i_address                             (nios2_qsys_0_instruction_master_address),                      //        instruction_master.address
		.i_read                                (nios2_qsys_0_instruction_master_read),                         //                          .read
		.i_readdata                            (nios2_qsys_0_instruction_master_readdata),                     //                          .readdata
		.i_waitrequest                         (nios2_qsys_0_instruction_master_waitrequest),                  //                          .waitrequest
		.d_irq                                 (nios2_qsys_0_d_irq_irq),                                       //                     d_irq.irq
		.jtag_debug_module_resetrequest        (nios2_qsys_0_jtag_debug_module_reset_reset),                   //   jtag_debug_module_reset.reset
		.jtag_debug_module_address             (mm_interconnect_0_nios2_qsys_0_jtag_debug_module_address),     //         jtag_debug_module.address
		.jtag_debug_module_byteenable          (mm_interconnect_0_nios2_qsys_0_jtag_debug_module_byteenable),  //                          .byteenable
		.jtag_debug_module_debugaccess         (mm_interconnect_0_nios2_qsys_0_jtag_debug_module_debugaccess), //                          .debugaccess
		.jtag_debug_module_read                (mm_interconnect_0_nios2_qsys_0_jtag_debug_module_read),        //                          .read
		.jtag_debug_module_readdata            (mm_interconnect_0_nios2_qsys_0_jtag_debug_module_readdata),    //                          .readdata
		.jtag_debug_module_waitrequest         (mm_interconnect_0_nios2_qsys_0_jtag_debug_module_waitrequest), //                          .waitrequest
		.jtag_debug_module_write               (mm_interconnect_0_nios2_qsys_0_jtag_debug_module_write),       //                          .write
		.jtag_debug_module_writedata           (mm_interconnect_0_nios2_qsys_0_jtag_debug_module_writedata),   //                          .writedata
		.no_ci_readra                          ()                                                              // custom_instruction_master.readra
	);

	nios_system_onchip_memory2_0 onchip_memory2_0 (
		.clk        (clk_clk),                                          //   clk1.clk
		.address    (mm_interconnect_0_onchip_memory2_0_s1_address),    //     s1.address
		.clken      (mm_interconnect_0_onchip_memory2_0_s1_clken),      //       .clken
		.chipselect (mm_interconnect_0_onchip_memory2_0_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_0_onchip_memory2_0_s1_write),      //       .write
		.readdata   (mm_interconnect_0_onchip_memory2_0_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_0_onchip_memory2_0_s1_writedata),  //       .writedata
		.byteenable (mm_interconnect_0_onchip_memory2_0_s1_byteenable), //       .byteenable
		.reset      (rst_controller_001_reset_out_reset),               // reset1.reset
		.reset_req  (rst_controller_001_reset_out_reset_req)            //       .reset_req
	);

	nios_system_otg_hpi_address otg_hpi_address (
		.clk        (clk_clk),                                         //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                 //               reset.reset_n
		.address    (mm_interconnect_0_otg_hpi_address_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_otg_hpi_address_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_otg_hpi_address_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_otg_hpi_address_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_otg_hpi_address_s1_readdata),   //                    .readdata
		.out_port   (otg_hpi_address_export)                           // external_connection.export
	);

	nios_system_otg_hpi_cs otg_hpi_cs (
		.clk        (clk_clk),                                    //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),            //               reset.reset_n
		.address    (mm_interconnect_0_otg_hpi_cs_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_otg_hpi_cs_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_otg_hpi_cs_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_otg_hpi_cs_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_otg_hpi_cs_s1_readdata),   //                    .readdata
		.out_port   (otg_hpi_cs_export)                           // external_connection.export
	);

	nios_system_otg_hpi_data otg_hpi_data (
		.clk        (clk_clk),                                      //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),              //               reset.reset_n
		.address    (mm_interconnect_0_otg_hpi_data_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_otg_hpi_data_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_otg_hpi_data_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_otg_hpi_data_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_otg_hpi_data_s1_readdata),   //                    .readdata
		.in_port    (otg_hpi_data_in_port),                         // external_connection.export
		.out_port   (otg_hpi_data_out_port)                         //                    .export
	);

	nios_system_otg_hpi_cs otg_hpi_r (
		.clk        (clk_clk),                                   //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),           //               reset.reset_n
		.address    (mm_interconnect_0_otg_hpi_r_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_otg_hpi_r_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_otg_hpi_r_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_otg_hpi_r_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_otg_hpi_r_s1_readdata),   //                    .readdata
		.out_port   (otg_hpi_r_export)                           // external_connection.export
	);

	nios_system_otg_hpi_cs otg_hpi_w (
		.clk        (clk_clk),                                   //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),           //               reset.reset_n
		.address    (mm_interconnect_0_otg_hpi_w_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_otg_hpi_w_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_otg_hpi_w_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_otg_hpi_w_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_otg_hpi_w_s1_readdata),   //                    .readdata
		.out_port   (otg_hpi_w_export)                           // external_connection.export
	);

	nios_system_EightBall poolcue (
		.clk        (clk_clk),                                 //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),         //               reset.reset_n
		.address    (mm_interconnect_0_poolcue_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_poolcue_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_poolcue_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_poolcue_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_poolcue_s1_readdata),   //                    .readdata
		.out_port   (poolcue_export)                           // external_connection.export
	);

	nios_system_sdram sdram (
		.clk            (sdram_pll_c0_clk),                         //   clk.clk
		.reset_n        (~rst_controller_002_reset_out_reset),      // reset.reset_n
		.az_addr        (mm_interconnect_0_sdram_s1_address),       //    s1.address
		.az_be_n        (~mm_interconnect_0_sdram_s1_byteenable),   //      .byteenable_n
		.az_cs          (mm_interconnect_0_sdram_s1_chipselect),    //      .chipselect
		.az_data        (mm_interconnect_0_sdram_s1_writedata),     //      .writedata
		.az_rd_n        (~mm_interconnect_0_sdram_s1_read),         //      .read_n
		.az_wr_n        (~mm_interconnect_0_sdram_s1_write),        //      .write_n
		.za_data        (mm_interconnect_0_sdram_s1_readdata),      //      .readdata
		.za_valid       (mm_interconnect_0_sdram_s1_readdatavalid), //      .readdatavalid
		.za_waitrequest (mm_interconnect_0_sdram_s1_waitrequest),   //      .waitrequest
		.zs_addr        (sdram_wire_addr),                          //  wire.export
		.zs_ba          (sdram_wire_ba),                            //      .export
		.zs_cas_n       (sdram_wire_cas_n),                         //      .export
		.zs_cke         (sdram_wire_cke),                           //      .export
		.zs_cs_n        (sdram_wire_cs_n),                          //      .export
		.zs_dq          (sdram_wire_dq),                            //      .export
		.zs_dqm         (sdram_wire_dqm),                           //      .export
		.zs_ras_n       (sdram_wire_ras_n),                         //      .export
		.zs_we_n        (sdram_wire_we_n)                           //      .export
	);

	nios_system_sdram_pll sdram_pll (
		.clk       (clk_clk),                                         //       inclk_interface.clk
		.reset     (rst_controller_001_reset_out_reset),              // inclk_interface_reset.reset
		.read      (mm_interconnect_0_sdram_pll_pll_slave_read),      //             pll_slave.read
		.write     (mm_interconnect_0_sdram_pll_pll_slave_write),     //                      .write
		.address   (mm_interconnect_0_sdram_pll_pll_slave_address),   //                      .address
		.readdata  (mm_interconnect_0_sdram_pll_pll_slave_readdata),  //                      .readdata
		.writedata (mm_interconnect_0_sdram_pll_pll_slave_writedata), //                      .writedata
		.c0        (sdram_pll_c0_clk),                                //                    c0.clk
		.c1        (sdram_clk_clk),                                   //                    c1.clk
		.areset    (),                                                //        areset_conduit.export
		.locked    (),                                                //        locked_conduit.export
		.phasedone ()                                                 //     phasedone_conduit.export
	);

	nios_system_sysid_qsys_0 sysid_qsys_0 (
		.clock    (clk_clk),                                               //           clk.clk
		.reset_n  (~rst_controller_001_reset_out_reset),                   //         reset.reset_n
		.readdata (mm_interconnect_0_sysid_qsys_0_control_slave_readdata), // control_slave.readdata
		.address  (mm_interconnect_0_sysid_qsys_0_control_slave_address)   //              .address
	);

	nios_system_reset reset (
		.clk      (clk_clk),                             //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),     //               reset.reset_n
		.address  (mm_interconnect_0_reset_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_reset_s1_readdata), //                    .readdata
		.in_port  (sys_reset_export)                     // external_connection.export
	);

	nios_system_reset hw_sig (
		.clk      (clk_clk),                              //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),      //               reset.reset_n
		.address  (mm_interconnect_0_hw_sig_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_hw_sig_s1_readdata), //                    .readdata
		.in_port  (hw_sig_export)                         // external_connection.export
	);

	nios_system_stick_direction stick_direction (
		.clk        (clk_clk),                                         //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                 //               reset.reset_n
		.address    (mm_interconnect_0_stick_direction_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_stick_direction_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_stick_direction_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_stick_direction_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_stick_direction_s1_readdata),   //                    .readdata
		.out_port   (stick_direction_export)                           // external_connection.export
	);

	nios_system_mm_interconnect_0 mm_interconnect_0 (
		.clk_0_clk_clk                                    (clk_clk),                                                      //                                  clk_0_clk.clk
		.sdram_pll_c0_clk                                 (sdram_pll_c0_clk),                                             //                               sdram_pll_c0.clk
		.jtag_uart_0_reset_reset_bridge_in_reset_reset    (rst_controller_reset_out_reset),                               //    jtag_uart_0_reset_reset_bridge_in_reset.reset
		.nios2_qsys_0_reset_n_reset_bridge_in_reset_reset (rst_controller_001_reset_out_reset),                           // nios2_qsys_0_reset_n_reset_bridge_in_reset.reset
		.sdram_reset_reset_bridge_in_reset_reset          (rst_controller_002_reset_out_reset),                           //          sdram_reset_reset_bridge_in_reset.reset
		.nios2_qsys_0_data_master_address                 (nios2_qsys_0_data_master_address),                             //                   nios2_qsys_0_data_master.address
		.nios2_qsys_0_data_master_waitrequest             (nios2_qsys_0_data_master_waitrequest),                         //                                           .waitrequest
		.nios2_qsys_0_data_master_byteenable              (nios2_qsys_0_data_master_byteenable),                          //                                           .byteenable
		.nios2_qsys_0_data_master_read                    (nios2_qsys_0_data_master_read),                                //                                           .read
		.nios2_qsys_0_data_master_readdata                (nios2_qsys_0_data_master_readdata),                            //                                           .readdata
		.nios2_qsys_0_data_master_write                   (nios2_qsys_0_data_master_write),                               //                                           .write
		.nios2_qsys_0_data_master_writedata               (nios2_qsys_0_data_master_writedata),                           //                                           .writedata
		.nios2_qsys_0_data_master_debugaccess             (nios2_qsys_0_data_master_debugaccess),                         //                                           .debugaccess
		.nios2_qsys_0_instruction_master_address          (nios2_qsys_0_instruction_master_address),                      //            nios2_qsys_0_instruction_master.address
		.nios2_qsys_0_instruction_master_waitrequest      (nios2_qsys_0_instruction_master_waitrequest),                  //                                           .waitrequest
		.nios2_qsys_0_instruction_master_read             (nios2_qsys_0_instruction_master_read),                         //                                           .read
		.nios2_qsys_0_instruction_master_readdata         (nios2_qsys_0_instruction_master_readdata),                     //                                           .readdata
		.cueBall_s1_address                               (mm_interconnect_0_cueball_s1_address),                         //                                 cueBall_s1.address
		.cueBall_s1_write                                 (mm_interconnect_0_cueball_s1_write),                           //                                           .write
		.cueBall_s1_readdata                              (mm_interconnect_0_cueball_s1_readdata),                        //                                           .readdata
		.cueBall_s1_writedata                             (mm_interconnect_0_cueball_s1_writedata),                       //                                           .writedata
		.cueBall_s1_chipselect                            (mm_interconnect_0_cueball_s1_chipselect),                      //                                           .chipselect
		.EightBall_s1_address                             (mm_interconnect_0_eightball_s1_address),                       //                               EightBall_s1.address
		.EightBall_s1_write                               (mm_interconnect_0_eightball_s1_write),                         //                                           .write
		.EightBall_s1_readdata                            (mm_interconnect_0_eightball_s1_readdata),                      //                                           .readdata
		.EightBall_s1_writedata                           (mm_interconnect_0_eightball_s1_writedata),                     //                                           .writedata
		.EightBall_s1_chipselect                          (mm_interconnect_0_eightball_s1_chipselect),                    //                                           .chipselect
		.ElevenBall_s1_address                            (mm_interconnect_0_elevenball_s1_address),                      //                              ElevenBall_s1.address
		.ElevenBall_s1_write                              (mm_interconnect_0_elevenball_s1_write),                        //                                           .write
		.ElevenBall_s1_readdata                           (mm_interconnect_0_elevenball_s1_readdata),                     //                                           .readdata
		.ElevenBall_s1_writedata                          (mm_interconnect_0_elevenball_s1_writedata),                    //                                           .writedata
		.ElevenBall_s1_chipselect                         (mm_interconnect_0_elevenball_s1_chipselect),                   //                                           .chipselect
		.FifteenBall_s1_address                           (mm_interconnect_0_fifteenball_s1_address),                     //                             FifteenBall_s1.address
		.FifteenBall_s1_write                             (mm_interconnect_0_fifteenball_s1_write),                       //                                           .write
		.FifteenBall_s1_readdata                          (mm_interconnect_0_fifteenball_s1_readdata),                    //                                           .readdata
		.FifteenBall_s1_writedata                         (mm_interconnect_0_fifteenball_s1_writedata),                   //                                           .writedata
		.FifteenBall_s1_chipselect                        (mm_interconnect_0_fifteenball_s1_chipselect),                  //                                           .chipselect
		.FiveBall_s1_address                              (mm_interconnect_0_fiveball_s1_address),                        //                                FiveBall_s1.address
		.FiveBall_s1_write                                (mm_interconnect_0_fiveball_s1_write),                          //                                           .write
		.FiveBall_s1_readdata                             (mm_interconnect_0_fiveball_s1_readdata),                       //                                           .readdata
		.FiveBall_s1_writedata                            (mm_interconnect_0_fiveball_s1_writedata),                      //                                           .writedata
		.FiveBall_s1_chipselect                           (mm_interconnect_0_fiveball_s1_chipselect),                     //                                           .chipselect
		.FourBall_s1_address                              (mm_interconnect_0_fourball_s1_address),                        //                                FourBall_s1.address
		.FourBall_s1_write                                (mm_interconnect_0_fourball_s1_write),                          //                                           .write
		.FourBall_s1_readdata                             (mm_interconnect_0_fourball_s1_readdata),                       //                                           .readdata
		.FourBall_s1_writedata                            (mm_interconnect_0_fourball_s1_writedata),                      //                                           .writedata
		.FourBall_s1_chipselect                           (mm_interconnect_0_fourball_s1_chipselect),                     //                                           .chipselect
		.FourteenBall_s1_address                          (mm_interconnect_0_fourteenball_s1_address),                    //                            FourteenBall_s1.address
		.FourteenBall_s1_write                            (mm_interconnect_0_fourteenball_s1_write),                      //                                           .write
		.FourteenBall_s1_readdata                         (mm_interconnect_0_fourteenball_s1_readdata),                   //                                           .readdata
		.FourteenBall_s1_writedata                        (mm_interconnect_0_fourteenball_s1_writedata),                  //                                           .writedata
		.FourteenBall_s1_chipselect                       (mm_interconnect_0_fourteenball_s1_chipselect),                 //                                           .chipselect
		.hw_sig_s1_address                                (mm_interconnect_0_hw_sig_s1_address),                          //                                  hw_sig_s1.address
		.hw_sig_s1_readdata                               (mm_interconnect_0_hw_sig_s1_readdata),                         //                                           .readdata
		.jtag_uart_0_avalon_jtag_slave_address            (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address),      //              jtag_uart_0_avalon_jtag_slave.address
		.jtag_uart_0_avalon_jtag_slave_write              (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write),        //                                           .write
		.jtag_uart_0_avalon_jtag_slave_read               (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read),         //                                           .read
		.jtag_uart_0_avalon_jtag_slave_readdata           (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata),     //                                           .readdata
		.jtag_uart_0_avalon_jtag_slave_writedata          (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata),    //                                           .writedata
		.jtag_uart_0_avalon_jtag_slave_waitrequest        (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest),  //                                           .waitrequest
		.jtag_uart_0_avalon_jtag_slave_chipselect         (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect),   //                                           .chipselect
		.keycode_s1_address                               (mm_interconnect_0_keycode_s1_address),                         //                                 keycode_s1.address
		.keycode_s1_write                                 (mm_interconnect_0_keycode_s1_write),                           //                                           .write
		.keycode_s1_readdata                              (mm_interconnect_0_keycode_s1_readdata),                        //                                           .readdata
		.keycode_s1_writedata                             (mm_interconnect_0_keycode_s1_writedata),                       //                                           .writedata
		.keycode_s1_chipselect                            (mm_interconnect_0_keycode_s1_chipselect),                      //                                           .chipselect
		.NineBall_s1_address                              (mm_interconnect_0_nineball_s1_address),                        //                                NineBall_s1.address
		.NineBall_s1_write                                (mm_interconnect_0_nineball_s1_write),                          //                                           .write
		.NineBall_s1_readdata                             (mm_interconnect_0_nineball_s1_readdata),                       //                                           .readdata
		.NineBall_s1_writedata                            (mm_interconnect_0_nineball_s1_writedata),                      //                                           .writedata
		.NineBall_s1_chipselect                           (mm_interconnect_0_nineball_s1_chipselect),                     //                                           .chipselect
		.nios2_qsys_0_jtag_debug_module_address           (mm_interconnect_0_nios2_qsys_0_jtag_debug_module_address),     //             nios2_qsys_0_jtag_debug_module.address
		.nios2_qsys_0_jtag_debug_module_write             (mm_interconnect_0_nios2_qsys_0_jtag_debug_module_write),       //                                           .write
		.nios2_qsys_0_jtag_debug_module_read              (mm_interconnect_0_nios2_qsys_0_jtag_debug_module_read),        //                                           .read
		.nios2_qsys_0_jtag_debug_module_readdata          (mm_interconnect_0_nios2_qsys_0_jtag_debug_module_readdata),    //                                           .readdata
		.nios2_qsys_0_jtag_debug_module_writedata         (mm_interconnect_0_nios2_qsys_0_jtag_debug_module_writedata),   //                                           .writedata
		.nios2_qsys_0_jtag_debug_module_byteenable        (mm_interconnect_0_nios2_qsys_0_jtag_debug_module_byteenable),  //                                           .byteenable
		.nios2_qsys_0_jtag_debug_module_waitrequest       (mm_interconnect_0_nios2_qsys_0_jtag_debug_module_waitrequest), //                                           .waitrequest
		.nios2_qsys_0_jtag_debug_module_debugaccess       (mm_interconnect_0_nios2_qsys_0_jtag_debug_module_debugaccess), //                                           .debugaccess
		.onchip_memory2_0_s1_address                      (mm_interconnect_0_onchip_memory2_0_s1_address),                //                        onchip_memory2_0_s1.address
		.onchip_memory2_0_s1_write                        (mm_interconnect_0_onchip_memory2_0_s1_write),                  //                                           .write
		.onchip_memory2_0_s1_readdata                     (mm_interconnect_0_onchip_memory2_0_s1_readdata),               //                                           .readdata
		.onchip_memory2_0_s1_writedata                    (mm_interconnect_0_onchip_memory2_0_s1_writedata),              //                                           .writedata
		.onchip_memory2_0_s1_byteenable                   (mm_interconnect_0_onchip_memory2_0_s1_byteenable),             //                                           .byteenable
		.onchip_memory2_0_s1_chipselect                   (mm_interconnect_0_onchip_memory2_0_s1_chipselect),             //                                           .chipselect
		.onchip_memory2_0_s1_clken                        (mm_interconnect_0_onchip_memory2_0_s1_clken),                  //                                           .clken
		.OneBall_s1_address                               (mm_interconnect_0_oneball_s1_address),                         //                                 OneBall_s1.address
		.OneBall_s1_write                                 (mm_interconnect_0_oneball_s1_write),                           //                                           .write
		.OneBall_s1_readdata                              (mm_interconnect_0_oneball_s1_readdata),                        //                                           .readdata
		.OneBall_s1_writedata                             (mm_interconnect_0_oneball_s1_writedata),                       //                                           .writedata
		.OneBall_s1_chipselect                            (mm_interconnect_0_oneball_s1_chipselect),                      //                                           .chipselect
		.otg_hpi_address_s1_address                       (mm_interconnect_0_otg_hpi_address_s1_address),                 //                         otg_hpi_address_s1.address
		.otg_hpi_address_s1_write                         (mm_interconnect_0_otg_hpi_address_s1_write),                   //                                           .write
		.otg_hpi_address_s1_readdata                      (mm_interconnect_0_otg_hpi_address_s1_readdata),                //                                           .readdata
		.otg_hpi_address_s1_writedata                     (mm_interconnect_0_otg_hpi_address_s1_writedata),               //                                           .writedata
		.otg_hpi_address_s1_chipselect                    (mm_interconnect_0_otg_hpi_address_s1_chipselect),              //                                           .chipselect
		.otg_hpi_cs_s1_address                            (mm_interconnect_0_otg_hpi_cs_s1_address),                      //                              otg_hpi_cs_s1.address
		.otg_hpi_cs_s1_write                              (mm_interconnect_0_otg_hpi_cs_s1_write),                        //                                           .write
		.otg_hpi_cs_s1_readdata                           (mm_interconnect_0_otg_hpi_cs_s1_readdata),                     //                                           .readdata
		.otg_hpi_cs_s1_writedata                          (mm_interconnect_0_otg_hpi_cs_s1_writedata),                    //                                           .writedata
		.otg_hpi_cs_s1_chipselect                         (mm_interconnect_0_otg_hpi_cs_s1_chipselect),                   //                                           .chipselect
		.otg_hpi_data_s1_address                          (mm_interconnect_0_otg_hpi_data_s1_address),                    //                            otg_hpi_data_s1.address
		.otg_hpi_data_s1_write                            (mm_interconnect_0_otg_hpi_data_s1_write),                      //                                           .write
		.otg_hpi_data_s1_readdata                         (mm_interconnect_0_otg_hpi_data_s1_readdata),                   //                                           .readdata
		.otg_hpi_data_s1_writedata                        (mm_interconnect_0_otg_hpi_data_s1_writedata),                  //                                           .writedata
		.otg_hpi_data_s1_chipselect                       (mm_interconnect_0_otg_hpi_data_s1_chipselect),                 //                                           .chipselect
		.otg_hpi_r_s1_address                             (mm_interconnect_0_otg_hpi_r_s1_address),                       //                               otg_hpi_r_s1.address
		.otg_hpi_r_s1_write                               (mm_interconnect_0_otg_hpi_r_s1_write),                         //                                           .write
		.otg_hpi_r_s1_readdata                            (mm_interconnect_0_otg_hpi_r_s1_readdata),                      //                                           .readdata
		.otg_hpi_r_s1_writedata                           (mm_interconnect_0_otg_hpi_r_s1_writedata),                     //                                           .writedata
		.otg_hpi_r_s1_chipselect                          (mm_interconnect_0_otg_hpi_r_s1_chipselect),                    //                                           .chipselect
		.otg_hpi_w_s1_address                             (mm_interconnect_0_otg_hpi_w_s1_address),                       //                               otg_hpi_w_s1.address
		.otg_hpi_w_s1_write                               (mm_interconnect_0_otg_hpi_w_s1_write),                         //                                           .write
		.otg_hpi_w_s1_readdata                            (mm_interconnect_0_otg_hpi_w_s1_readdata),                      //                                           .readdata
		.otg_hpi_w_s1_writedata                           (mm_interconnect_0_otg_hpi_w_s1_writedata),                     //                                           .writedata
		.otg_hpi_w_s1_chipselect                          (mm_interconnect_0_otg_hpi_w_s1_chipselect),                    //                                           .chipselect
		.poolcue_s1_address                               (mm_interconnect_0_poolcue_s1_address),                         //                                 poolcue_s1.address
		.poolcue_s1_write                                 (mm_interconnect_0_poolcue_s1_write),                           //                                           .write
		.poolcue_s1_readdata                              (mm_interconnect_0_poolcue_s1_readdata),                        //                                           .readdata
		.poolcue_s1_writedata                             (mm_interconnect_0_poolcue_s1_writedata),                       //                                           .writedata
		.poolcue_s1_chipselect                            (mm_interconnect_0_poolcue_s1_chipselect),                      //                                           .chipselect
		.reset_s1_address                                 (mm_interconnect_0_reset_s1_address),                           //                                   reset_s1.address
		.reset_s1_readdata                                (mm_interconnect_0_reset_s1_readdata),                          //                                           .readdata
		.sdram_s1_address                                 (mm_interconnect_0_sdram_s1_address),                           //                                   sdram_s1.address
		.sdram_s1_write                                   (mm_interconnect_0_sdram_s1_write),                             //                                           .write
		.sdram_s1_read                                    (mm_interconnect_0_sdram_s1_read),                              //                                           .read
		.sdram_s1_readdata                                (mm_interconnect_0_sdram_s1_readdata),                          //                                           .readdata
		.sdram_s1_writedata                               (mm_interconnect_0_sdram_s1_writedata),                         //                                           .writedata
		.sdram_s1_byteenable                              (mm_interconnect_0_sdram_s1_byteenable),                        //                                           .byteenable
		.sdram_s1_readdatavalid                           (mm_interconnect_0_sdram_s1_readdatavalid),                     //                                           .readdatavalid
		.sdram_s1_waitrequest                             (mm_interconnect_0_sdram_s1_waitrequest),                       //                                           .waitrequest
		.sdram_s1_chipselect                              (mm_interconnect_0_sdram_s1_chipselect),                        //                                           .chipselect
		.sdram_pll_pll_slave_address                      (mm_interconnect_0_sdram_pll_pll_slave_address),                //                        sdram_pll_pll_slave.address
		.sdram_pll_pll_slave_write                        (mm_interconnect_0_sdram_pll_pll_slave_write),                  //                                           .write
		.sdram_pll_pll_slave_read                         (mm_interconnect_0_sdram_pll_pll_slave_read),                   //                                           .read
		.sdram_pll_pll_slave_readdata                     (mm_interconnect_0_sdram_pll_pll_slave_readdata),               //                                           .readdata
		.sdram_pll_pll_slave_writedata                    (mm_interconnect_0_sdram_pll_pll_slave_writedata),              //                                           .writedata
		.SevenBall_s1_address                             (mm_interconnect_0_sevenball_s1_address),                       //                               SevenBall_s1.address
		.SevenBall_s1_write                               (mm_interconnect_0_sevenball_s1_write),                         //                                           .write
		.SevenBall_s1_readdata                            (mm_interconnect_0_sevenball_s1_readdata),                      //                                           .readdata
		.SevenBall_s1_writedata                           (mm_interconnect_0_sevenball_s1_writedata),                     //                                           .writedata
		.SevenBall_s1_chipselect                          (mm_interconnect_0_sevenball_s1_chipselect),                    //                                           .chipselect
		.SixBall_s1_address                               (mm_interconnect_0_sixball_s1_address),                         //                                 SixBall_s1.address
		.SixBall_s1_write                                 (mm_interconnect_0_sixball_s1_write),                           //                                           .write
		.SixBall_s1_readdata                              (mm_interconnect_0_sixball_s1_readdata),                        //                                           .readdata
		.SixBall_s1_writedata                             (mm_interconnect_0_sixball_s1_writedata),                       //                                           .writedata
		.SixBall_s1_chipselect                            (mm_interconnect_0_sixball_s1_chipselect),                      //                                           .chipselect
		.stick_direction_s1_address                       (mm_interconnect_0_stick_direction_s1_address),                 //                         stick_direction_s1.address
		.stick_direction_s1_write                         (mm_interconnect_0_stick_direction_s1_write),                   //                                           .write
		.stick_direction_s1_readdata                      (mm_interconnect_0_stick_direction_s1_readdata),                //                                           .readdata
		.stick_direction_s1_writedata                     (mm_interconnect_0_stick_direction_s1_writedata),               //                                           .writedata
		.stick_direction_s1_chipselect                    (mm_interconnect_0_stick_direction_s1_chipselect),              //                                           .chipselect
		.sysid_qsys_0_control_slave_address               (mm_interconnect_0_sysid_qsys_0_control_slave_address),         //                 sysid_qsys_0_control_slave.address
		.sysid_qsys_0_control_slave_readdata              (mm_interconnect_0_sysid_qsys_0_control_slave_readdata),        //                                           .readdata
		.TenBall_s1_address                               (mm_interconnect_0_tenball_s1_address),                         //                                 TenBall_s1.address
		.TenBall_s1_write                                 (mm_interconnect_0_tenball_s1_write),                           //                                           .write
		.TenBall_s1_readdata                              (mm_interconnect_0_tenball_s1_readdata),                        //                                           .readdata
		.TenBall_s1_writedata                             (mm_interconnect_0_tenball_s1_writedata),                       //                                           .writedata
		.TenBall_s1_chipselect                            (mm_interconnect_0_tenball_s1_chipselect),                      //                                           .chipselect
		.ThirteenBall_s1_address                          (mm_interconnect_0_thirteenball_s1_address),                    //                            ThirteenBall_s1.address
		.ThirteenBall_s1_write                            (mm_interconnect_0_thirteenball_s1_write),                      //                                           .write
		.ThirteenBall_s1_readdata                         (mm_interconnect_0_thirteenball_s1_readdata),                   //                                           .readdata
		.ThirteenBall_s1_writedata                        (mm_interconnect_0_thirteenball_s1_writedata),                  //                                           .writedata
		.ThirteenBall_s1_chipselect                       (mm_interconnect_0_thirteenball_s1_chipselect),                 //                                           .chipselect
		.ThreeBall_s1_address                             (mm_interconnect_0_threeball_s1_address),                       //                               ThreeBall_s1.address
		.ThreeBall_s1_write                               (mm_interconnect_0_threeball_s1_write),                         //                                           .write
		.ThreeBall_s1_readdata                            (mm_interconnect_0_threeball_s1_readdata),                      //                                           .readdata
		.ThreeBall_s1_writedata                           (mm_interconnect_0_threeball_s1_writedata),                     //                                           .writedata
		.ThreeBall_s1_chipselect                          (mm_interconnect_0_threeball_s1_chipselect),                    //                                           .chipselect
		.TwelveBall_s1_address                            (mm_interconnect_0_twelveball_s1_address),                      //                              TwelveBall_s1.address
		.TwelveBall_s1_write                              (mm_interconnect_0_twelveball_s1_write),                        //                                           .write
		.TwelveBall_s1_readdata                           (mm_interconnect_0_twelveball_s1_readdata),                     //                                           .readdata
		.TwelveBall_s1_writedata                          (mm_interconnect_0_twelveball_s1_writedata),                    //                                           .writedata
		.TwelveBall_s1_chipselect                         (mm_interconnect_0_twelveball_s1_chipselect),                   //                                           .chipselect
		.TwoBall_s1_address                               (mm_interconnect_0_twoball_s1_address),                         //                                 TwoBall_s1.address
		.TwoBall_s1_write                                 (mm_interconnect_0_twoball_s1_write),                           //                                           .write
		.TwoBall_s1_readdata                              (mm_interconnect_0_twoball_s1_readdata),                        //                                           .readdata
		.TwoBall_s1_writedata                             (mm_interconnect_0_twoball_s1_writedata),                       //                                           .writedata
		.TwoBall_s1_chipselect                            (mm_interconnect_0_twoball_s1_chipselect)                       //                                           .chipselect
	);

	nios_system_irq_mapper irq_mapper (
		.clk           (clk_clk),                            //       clk.clk
		.reset         (rst_controller_001_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),           // receiver0.irq
		.sender_irq    (nios2_qsys_0_d_irq_irq)              //    sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                             // reset_in0.reset
		.reset_in1      (nios2_qsys_0_jtag_debug_module_reset_reset), // reset_in1.reset
		.clk            (clk_clk),                                    //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),             // reset_out.reset
		.reset_req      (),                                           // (terminated)
		.reset_req_in0  (1'b0),                                       // (terminated)
		.reset_req_in1  (1'b0),                                       // (terminated)
		.reset_in2      (1'b0),                                       // (terminated)
		.reset_req_in2  (1'b0),                                       // (terminated)
		.reset_in3      (1'b0),                                       // (terminated)
		.reset_req_in3  (1'b0),                                       // (terminated)
		.reset_in4      (1'b0),                                       // (terminated)
		.reset_req_in4  (1'b0),                                       // (terminated)
		.reset_in5      (1'b0),                                       // (terminated)
		.reset_req_in5  (1'b0),                                       // (terminated)
		.reset_in6      (1'b0),                                       // (terminated)
		.reset_req_in6  (1'b0),                                       // (terminated)
		.reset_in7      (1'b0),                                       // (terminated)
		.reset_req_in7  (1'b0),                                       // (terminated)
		.reset_in8      (1'b0),                                       // (terminated)
		.reset_req_in8  (1'b0),                                       // (terminated)
		.reset_in9      (1'b0),                                       // (terminated)
		.reset_req_in9  (1'b0),                                       // (terminated)
		.reset_in10     (1'b0),                                       // (terminated)
		.reset_req_in10 (1'b0),                                       // (terminated)
		.reset_in11     (1'b0),                                       // (terminated)
		.reset_req_in11 (1'b0),                                       // (terminated)
		.reset_in12     (1'b0),                                       // (terminated)
		.reset_req_in12 (1'b0),                                       // (terminated)
		.reset_in13     (1'b0),                                       // (terminated)
		.reset_req_in13 (1'b0),                                       // (terminated)
		.reset_in14     (1'b0),                                       // (terminated)
		.reset_req_in14 (1'b0),                                       // (terminated)
		.reset_in15     (1'b0),                                       // (terminated)
		.reset_req_in15 (1'b0)                                        // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_001 (
		.reset_in0      (~reset_reset_n),                         // reset_in0.reset
		.clk            (clk_clk),                                //       clk.clk
		.reset_out      (rst_controller_001_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_001_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                                   // (terminated)
		.reset_in1      (1'b0),                                   // (terminated)
		.reset_req_in1  (1'b0),                                   // (terminated)
		.reset_in2      (1'b0),                                   // (terminated)
		.reset_req_in2  (1'b0),                                   // (terminated)
		.reset_in3      (1'b0),                                   // (terminated)
		.reset_req_in3  (1'b0),                                   // (terminated)
		.reset_in4      (1'b0),                                   // (terminated)
		.reset_req_in4  (1'b0),                                   // (terminated)
		.reset_in5      (1'b0),                                   // (terminated)
		.reset_req_in5  (1'b0),                                   // (terminated)
		.reset_in6      (1'b0),                                   // (terminated)
		.reset_req_in6  (1'b0),                                   // (terminated)
		.reset_in7      (1'b0),                                   // (terminated)
		.reset_req_in7  (1'b0),                                   // (terminated)
		.reset_in8      (1'b0),                                   // (terminated)
		.reset_req_in8  (1'b0),                                   // (terminated)
		.reset_in9      (1'b0),                                   // (terminated)
		.reset_req_in9  (1'b0),                                   // (terminated)
		.reset_in10     (1'b0),                                   // (terminated)
		.reset_req_in10 (1'b0),                                   // (terminated)
		.reset_in11     (1'b0),                                   // (terminated)
		.reset_req_in11 (1'b0),                                   // (terminated)
		.reset_in12     (1'b0),                                   // (terminated)
		.reset_req_in12 (1'b0),                                   // (terminated)
		.reset_in13     (1'b0),                                   // (terminated)
		.reset_req_in13 (1'b0),                                   // (terminated)
		.reset_in14     (1'b0),                                   // (terminated)
		.reset_req_in14 (1'b0),                                   // (terminated)
		.reset_in15     (1'b0),                                   // (terminated)
		.reset_req_in15 (1'b0)                                    // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_002 (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.clk            (sdram_pll_c0_clk),                   //       clk.clk
		.reset_out      (rst_controller_002_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

endmodule
