library verilog;
use verilog.vl_types.all;
entity nios_system_mm_interconnect_0 is
    port(
        clk_0_clk_clk   : in     vl_logic;
        sdram_pll_c0_clk: in     vl_logic;
        jtag_uart_0_reset_reset_bridge_in_reset_reset: in     vl_logic;
        nios2_qsys_0_reset_n_reset_bridge_in_reset_reset: in     vl_logic;
        sdram_reset_reset_bridge_in_reset_reset: in     vl_logic;
        nios2_qsys_0_data_master_address: in     vl_logic_vector(28 downto 0);
        nios2_qsys_0_data_master_waitrequest: out    vl_logic;
        nios2_qsys_0_data_master_byteenable: in     vl_logic_vector(3 downto 0);
        nios2_qsys_0_data_master_read: in     vl_logic;
        nios2_qsys_0_data_master_readdata: out    vl_logic_vector(31 downto 0);
        nios2_qsys_0_data_master_write: in     vl_logic;
        nios2_qsys_0_data_master_writedata: in     vl_logic_vector(31 downto 0);
        nios2_qsys_0_data_master_debugaccess: in     vl_logic;
        nios2_qsys_0_instruction_master_address: in     vl_logic_vector(28 downto 0);
        nios2_qsys_0_instruction_master_waitrequest: out    vl_logic;
        nios2_qsys_0_instruction_master_read: in     vl_logic;
        nios2_qsys_0_instruction_master_readdata: out    vl_logic_vector(31 downto 0);
        cueBall_s1_address: out    vl_logic_vector(1 downto 0);
        cueBall_s1_write: out    vl_logic;
        cueBall_s1_readdata: in     vl_logic_vector(31 downto 0);
        cueBall_s1_writedata: out    vl_logic_vector(31 downto 0);
        cueBall_s1_chipselect: out    vl_logic;
        EightBall_s1_address: out    vl_logic_vector(1 downto 0);
        EightBall_s1_write: out    vl_logic;
        EightBall_s1_readdata: in     vl_logic_vector(31 downto 0);
        EightBall_s1_writedata: out    vl_logic_vector(31 downto 0);
        EightBall_s1_chipselect: out    vl_logic;
        ElevenBall_s1_address: out    vl_logic_vector(1 downto 0);
        ElevenBall_s1_write: out    vl_logic;
        ElevenBall_s1_readdata: in     vl_logic_vector(31 downto 0);
        ElevenBall_s1_writedata: out    vl_logic_vector(31 downto 0);
        ElevenBall_s1_chipselect: out    vl_logic;
        FifteenBall_s1_address: out    vl_logic_vector(1 downto 0);
        FifteenBall_s1_write: out    vl_logic;
        FifteenBall_s1_readdata: in     vl_logic_vector(31 downto 0);
        FifteenBall_s1_writedata: out    vl_logic_vector(31 downto 0);
        FifteenBall_s1_chipselect: out    vl_logic;
        FiveBall_s1_address: out    vl_logic_vector(1 downto 0);
        FiveBall_s1_write: out    vl_logic;
        FiveBall_s1_readdata: in     vl_logic_vector(31 downto 0);
        FiveBall_s1_writedata: out    vl_logic_vector(31 downto 0);
        FiveBall_s1_chipselect: out    vl_logic;
        FourBall_s1_address: out    vl_logic_vector(1 downto 0);
        FourBall_s1_write: out    vl_logic;
        FourBall_s1_readdata: in     vl_logic_vector(31 downto 0);
        FourBall_s1_writedata: out    vl_logic_vector(31 downto 0);
        FourBall_s1_chipselect: out    vl_logic;
        FourteenBall_s1_address: out    vl_logic_vector(1 downto 0);
        FourteenBall_s1_write: out    vl_logic;
        FourteenBall_s1_readdata: in     vl_logic_vector(31 downto 0);
        FourteenBall_s1_writedata: out    vl_logic_vector(31 downto 0);
        FourteenBall_s1_chipselect: out    vl_logic;
        hw_sig_s1_address: out    vl_logic_vector(1 downto 0);
        hw_sig_s1_readdata: in     vl_logic_vector(31 downto 0);
        jtag_uart_0_avalon_jtag_slave_address: out    vl_logic_vector(0 downto 0);
        jtag_uart_0_avalon_jtag_slave_write: out    vl_logic;
        jtag_uart_0_avalon_jtag_slave_read: out    vl_logic;
        jtag_uart_0_avalon_jtag_slave_readdata: in     vl_logic_vector(31 downto 0);
        jtag_uart_0_avalon_jtag_slave_writedata: out    vl_logic_vector(31 downto 0);
        jtag_uart_0_avalon_jtag_slave_waitrequest: in     vl_logic;
        jtag_uart_0_avalon_jtag_slave_chipselect: out    vl_logic;
        keycode_s1_address: out    vl_logic_vector(1 downto 0);
        keycode_s1_write: out    vl_logic;
        keycode_s1_readdata: in     vl_logic_vector(31 downto 0);
        keycode_s1_writedata: out    vl_logic_vector(31 downto 0);
        keycode_s1_chipselect: out    vl_logic;
        NineBall_s1_address: out    vl_logic_vector(1 downto 0);
        NineBall_s1_write: out    vl_logic;
        NineBall_s1_readdata: in     vl_logic_vector(31 downto 0);
        NineBall_s1_writedata: out    vl_logic_vector(31 downto 0);
        NineBall_s1_chipselect: out    vl_logic;
        nios2_qsys_0_jtag_debug_module_address: out    vl_logic_vector(8 downto 0);
        nios2_qsys_0_jtag_debug_module_write: out    vl_logic;
        nios2_qsys_0_jtag_debug_module_read: out    vl_logic;
        nios2_qsys_0_jtag_debug_module_readdata: in     vl_logic_vector(31 downto 0);
        nios2_qsys_0_jtag_debug_module_writedata: out    vl_logic_vector(31 downto 0);
        nios2_qsys_0_jtag_debug_module_byteenable: out    vl_logic_vector(3 downto 0);
        nios2_qsys_0_jtag_debug_module_waitrequest: in     vl_logic;
        nios2_qsys_0_jtag_debug_module_debugaccess: out    vl_logic;
        onchip_memory2_0_s1_address: out    vl_logic_vector(1 downto 0);
        onchip_memory2_0_s1_write: out    vl_logic;
        onchip_memory2_0_s1_readdata: in     vl_logic_vector(31 downto 0);
        onchip_memory2_0_s1_writedata: out    vl_logic_vector(31 downto 0);
        onchip_memory2_0_s1_byteenable: out    vl_logic_vector(3 downto 0);
        onchip_memory2_0_s1_chipselect: out    vl_logic;
        onchip_memory2_0_s1_clken: out    vl_logic;
        OneBall_s1_address: out    vl_logic_vector(1 downto 0);
        OneBall_s1_write: out    vl_logic;
        OneBall_s1_readdata: in     vl_logic_vector(31 downto 0);
        OneBall_s1_writedata: out    vl_logic_vector(31 downto 0);
        OneBall_s1_chipselect: out    vl_logic;
        otg_hpi_address_s1_address: out    vl_logic_vector(1 downto 0);
        otg_hpi_address_s1_write: out    vl_logic;
        otg_hpi_address_s1_readdata: in     vl_logic_vector(31 downto 0);
        otg_hpi_address_s1_writedata: out    vl_logic_vector(31 downto 0);
        otg_hpi_address_s1_chipselect: out    vl_logic;
        otg_hpi_cs_s1_address: out    vl_logic_vector(1 downto 0);
        otg_hpi_cs_s1_write: out    vl_logic;
        otg_hpi_cs_s1_readdata: in     vl_logic_vector(31 downto 0);
        otg_hpi_cs_s1_writedata: out    vl_logic_vector(31 downto 0);
        otg_hpi_cs_s1_chipselect: out    vl_logic;
        otg_hpi_data_s1_address: out    vl_logic_vector(1 downto 0);
        otg_hpi_data_s1_write: out    vl_logic;
        otg_hpi_data_s1_readdata: in     vl_logic_vector(31 downto 0);
        otg_hpi_data_s1_writedata: out    vl_logic_vector(31 downto 0);
        otg_hpi_data_s1_chipselect: out    vl_logic;
        otg_hpi_r_s1_address: out    vl_logic_vector(1 downto 0);
        otg_hpi_r_s1_write: out    vl_logic;
        otg_hpi_r_s1_readdata: in     vl_logic_vector(31 downto 0);
        otg_hpi_r_s1_writedata: out    vl_logic_vector(31 downto 0);
        otg_hpi_r_s1_chipselect: out    vl_logic;
        otg_hpi_w_s1_address: out    vl_logic_vector(1 downto 0);
        otg_hpi_w_s1_write: out    vl_logic;
        otg_hpi_w_s1_readdata: in     vl_logic_vector(31 downto 0);
        otg_hpi_w_s1_writedata: out    vl_logic_vector(31 downto 0);
        otg_hpi_w_s1_chipselect: out    vl_logic;
        poolcue_s1_address: out    vl_logic_vector(1 downto 0);
        poolcue_s1_write: out    vl_logic;
        poolcue_s1_readdata: in     vl_logic_vector(31 downto 0);
        poolcue_s1_writedata: out    vl_logic_vector(31 downto 0);
        poolcue_s1_chipselect: out    vl_logic;
        reset_s1_address: out    vl_logic_vector(1 downto 0);
        reset_s1_readdata: in     vl_logic_vector(31 downto 0);
        sdram_s1_address: out    vl_logic_vector(24 downto 0);
        sdram_s1_write  : out    vl_logic;
        sdram_s1_read   : out    vl_logic;
        sdram_s1_readdata: in     vl_logic_vector(31 downto 0);
        sdram_s1_writedata: out    vl_logic_vector(31 downto 0);
        sdram_s1_byteenable: out    vl_logic_vector(3 downto 0);
        sdram_s1_readdatavalid: in     vl_logic;
        sdram_s1_waitrequest: in     vl_logic;
        sdram_s1_chipselect: out    vl_logic;
        sdram_pll_pll_slave_address: out    vl_logic_vector(1 downto 0);
        sdram_pll_pll_slave_write: out    vl_logic;
        sdram_pll_pll_slave_read: out    vl_logic;
        sdram_pll_pll_slave_readdata: in     vl_logic_vector(31 downto 0);
        sdram_pll_pll_slave_writedata: out    vl_logic_vector(31 downto 0);
        SevenBall_s1_address: out    vl_logic_vector(1 downto 0);
        SevenBall_s1_write: out    vl_logic;
        SevenBall_s1_readdata: in     vl_logic_vector(31 downto 0);
        SevenBall_s1_writedata: out    vl_logic_vector(31 downto 0);
        SevenBall_s1_chipselect: out    vl_logic;
        SixBall_s1_address: out    vl_logic_vector(1 downto 0);
        SixBall_s1_write: out    vl_logic;
        SixBall_s1_readdata: in     vl_logic_vector(31 downto 0);
        SixBall_s1_writedata: out    vl_logic_vector(31 downto 0);
        SixBall_s1_chipselect: out    vl_logic;
        stick_direction_s1_address: out    vl_logic_vector(1 downto 0);
        stick_direction_s1_write: out    vl_logic;
        stick_direction_s1_readdata: in     vl_logic_vector(31 downto 0);
        stick_direction_s1_writedata: out    vl_logic_vector(31 downto 0);
        stick_direction_s1_chipselect: out    vl_logic;
        sysid_qsys_0_control_slave_address: out    vl_logic_vector(0 downto 0);
        sysid_qsys_0_control_slave_readdata: in     vl_logic_vector(31 downto 0);
        TenBall_s1_address: out    vl_logic_vector(1 downto 0);
        TenBall_s1_write: out    vl_logic;
        TenBall_s1_readdata: in     vl_logic_vector(31 downto 0);
        TenBall_s1_writedata: out    vl_logic_vector(31 downto 0);
        TenBall_s1_chipselect: out    vl_logic;
        ThirteenBall_s1_address: out    vl_logic_vector(1 downto 0);
        ThirteenBall_s1_write: out    vl_logic;
        ThirteenBall_s1_readdata: in     vl_logic_vector(31 downto 0);
        ThirteenBall_s1_writedata: out    vl_logic_vector(31 downto 0);
        ThirteenBall_s1_chipselect: out    vl_logic;
        ThreeBall_s1_address: out    vl_logic_vector(1 downto 0);
        ThreeBall_s1_write: out    vl_logic;
        ThreeBall_s1_readdata: in     vl_logic_vector(31 downto 0);
        ThreeBall_s1_writedata: out    vl_logic_vector(31 downto 0);
        ThreeBall_s1_chipselect: out    vl_logic;
        TwelveBall_s1_address: out    vl_logic_vector(1 downto 0);
        TwelveBall_s1_write: out    vl_logic;
        TwelveBall_s1_readdata: in     vl_logic_vector(31 downto 0);
        TwelveBall_s1_writedata: out    vl_logic_vector(31 downto 0);
        TwelveBall_s1_chipselect: out    vl_logic;
        TwoBall_s1_address: out    vl_logic_vector(1 downto 0);
        TwoBall_s1_write: out    vl_logic;
        TwoBall_s1_readdata: in     vl_logic_vector(31 downto 0);
        TwoBall_s1_writedata: out    vl_logic_vector(31 downto 0);
        TwoBall_s1_chipselect: out    vl_logic
    );
end nios_system_mm_interconnect_0;
